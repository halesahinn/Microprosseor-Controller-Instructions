module control(in,regdest,alusrc,memtoreg,regwrite,memread,memwrite,branch,ext,jump,jspa,aluop1,aluop2);
input [5:0] in;
output regdest,alusrc,memtoreg,regwrite,memread,memwrite,branch,ext,jump,jspa,aluop1,aluop2;
wire rformat,lw,sw,beq,bgez,xori,brn;
assign rformat=~|in;
assign lw=in[5]& (~in[4])&(~in[3])&(~in[2])&in[1]&in[0];
assign sw=in[5]& (~in[4])&in[3]&(~in[2])&in[1]&in[0];
assign beq=~in[5]& (~in[4])&(~in[3])&in[2]&(~in[1])&(~in[0]);
assign bgez=in[5]& (~in[4])&(~in[3])&in[2]&(in[1])&(in[0]);
assign xori=~in[5]& (~in[4])&(in[3])&in[2]&(in[1])&(~in[0]);
assign balz=~in[5]& (in[4])&(in[3])&~(in[2])&(in[1])&(~in[0]);
assign jspal=~in[5]& (in[4])&~(in[3])&~(in[2])&(in[1])&(in[0]);
assign regdest=rformat;
assign alusrc=lw|sw|xori;
assign memtoreg=lw;
assign regwrite=rformat|lw|xori;
assign memread=lw|jspal;
assign memwrite=sw|jspal;
assign branch=beq|bgez|brn;
assign ext=xori;
assign jspa=jspal;
assign jump=balz|jspal;
assign aluop1=rformat|xori;
assign aluop2=beq|bgez|xori|balz;
endmodule
